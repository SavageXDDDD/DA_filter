module main ();




endmodule