`define FIRST_SUBFILTER
`define LAST_SUBFILTER